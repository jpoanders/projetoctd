-- Teste
